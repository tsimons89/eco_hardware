`include "eco_includes.svh"

module eco_features_tb;

   eco_features my_eco_features(.*);

   task read_adaboost_file();
      
   endtask
endmodule
