module tree();

endmodule
