`ifndef ECO_INCLUDES
 `define ECO_INCLUDES
 `include "globals.svh"
 `include "eco_types.sv"
 `include "x_shift.sv"
 `include "y_shift.sv"
 `include "features.sv"
 `include "tree_node_data.sv"
 `include "tree_structure.sv"
 `include "tree_prediction_data.sv"
 `include "tree_node_compare.sv"
 `include "tree.sv"
 `include "tree_node.sv"
 `include "forest.sv"
 `include "forest_prediction.sv"
 `include "features_selection.sv"
 `include "ada_boost.sv"
`endif
