module eco_features(input clk,rst,px_stobe,load_node,load_prediction,set_feature_index,
		[`PIXEL_WIDTH - 1:0] px_value,[`FEATURE_INDEX_WIDTH] feature_index,
		node_data node_in,
		[`PREDICTION_WIDTH - 1:0] prediction_in,
		[`TREE_NUM_WIDTH - 1:0] tree_num,[`FOREST_NUM_WIDTH - 1:0] forest_num
		);
endmodule
